module jk_ff(input clk, j, k, output reg q);
    always @(posedge clk) begin
        case({j,k})
            2'b00: q <= q;
            2'b01: q <= 0;
            2'b10: q <= 1;
            2'b11: q <= ~q;
        endcase
    end
endmodule

module sr_ff(input clk, s, r, output reg q);
    always @(posedge clk) begin
        if (s & ~r) q <= 1;
        else if (~s & r) q <= 0;
        else if (s & r) q <= 1'bx;
    end
endmodule
