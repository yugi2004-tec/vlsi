module d_ff_en(input clk, en, d, output reg q);
    always @(posedge clk) begin
        if (en)
            q <= d;
    end
endmodule
